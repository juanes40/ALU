library verilog;
use verilog.vl_types.all;
entity alufinal_vlg_vec_tst is
end alufinal_vlg_vec_tst;
